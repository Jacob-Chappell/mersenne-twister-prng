module test();

endmodule
